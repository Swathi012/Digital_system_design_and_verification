module or_gate(input bit a, input bit b, output bit c);
assign c = a | b;
endmodule
