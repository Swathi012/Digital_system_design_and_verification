module not_gate(input bit a, output bit not_a);
assign not_a = ~a;
endmodule;

